`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Aleksander Kaminski
// 
// Create Date:    04:23:50 07/08/2014 
// Design Name:		Braindfuck CPU
// Module Name:    brainfuck_cpu_tb 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module brainfuck_cpu_tb();

	reg clk;
	reg rst;
	wire [7:0] data_i;
	wire [7:0] data_o;
	reg [2:0] rom_i;
	wire [10:0] data_addr_o;
	wire [6:0] rom_addr_o;
	wire rd;
	wire wr;
	wire mreq;
	wire ioreq;
	reg ready;

	reg ready_fsm, ready_fsm_next;

	brainfuck_cpu #(11,7,8) uut(clk, rst, data_i, data_o, rom_i, data_addr_o, rom_addr_o, rd, wr, mreq, ioreq, ready);

	always @(posedge clk, posedge rst) begin
		if (rst)
			ready_fsm <= 0;
		else
			ready_fsm <= ready_fsm_next;
	end

	always @(*) begin
		case (ready_fsm)
			0: begin
					ready <= 0;
					if (rd||wr)
						ready_fsm_next <= 1;
					else
						ready_fsm_next <= 0;
				end
			1: begin
					ready <= 1;
					ready_fsm_next <= 0;
				end
		endcase
	end

	initial begin
		rst <= 1'b1;
		clk <= 1'b0;
		#100 rst <= 1'b0;
	end

	always
		#1 clk <= ~clk;

	RAMB16_S9 #(
      .INIT(9'h000),  // Value of output RAM registers at startup
      .SRVAL(9'h000), // Output value upon SSR assertion
      .WRITE_MODE("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE

      // The forllowing INIT_xx declarations specify the initial contents of the RAM
      // Address 0 to 511
      .INIT_00(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_01(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_02(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_03(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_04(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_05(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_06(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_07(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_08(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_09(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_0A(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_0B(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_0C(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_0D(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_0E(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_0F(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      // Address 512 to 1023
      .INIT_10(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_11(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_12(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_13(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_14(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_15(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_16(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_17(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_18(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_19(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_1A(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_1B(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_1C(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_1D(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_1E(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_1F(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      // Address 1024 to 1535
      .INIT_20(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_21(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_22(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_23(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_24(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_25(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_26(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_27(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_28(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_29(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_2A(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_2B(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_2C(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_2D(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_2E(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_2F(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      // Address 1536 to 2047
      .INIT_30(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_31(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_32(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_33(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_34(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_35(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_36(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_37(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_38(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_39(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_3A(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_3B(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_3C(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_3D(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_3E(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_3F(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),

      // The next set of INITP_xx are for the parity bits
      // Address 0 to 511
      .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 512 to 1023
      .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 1024 to 1535
      .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 1536 to 2047
      .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000)
   ) RAMB16_S9_inst (
      .DO(data_i),      // 8-bit Data Output
      .DOP(),    // 1-bit parity Output
      .ADDR(data_addr_o),  // 11-bit Address Input
      .CLK(clk),    // Clock
      .DI(data_o),      // 8-bit Data Input
      .DIP(1'b0),    // 1-bit parity Input
      .EN(mreq),      // RAM Enable Input
      .SSR(rst),    // Synchronous Set/Reset Input
      .WE(wr)       // Write Enable Input
   );

	always @(negedge clk)
		if (wr && ioreq)
			$display("%c", data_o);

	always @(*) begin
		case (rom_addr_o)
			7'd0: rom_i <= 3'b010;    //+
			7'd1: rom_i <= 3'b010;    //+
			7'd2: rom_i <= 3'b010;    //+
			7'd3: rom_i <= 3'b010;    //+
			7'd4: rom_i <= 3'b010;    //+
			7'd5: rom_i <= 3'b010;    //+
			7'd6: rom_i <= 3'b010;    //+
			7'd7: rom_i <= 3'b010;    //+
			7'd8: rom_i <= 3'b010;    //+
			7'd9: rom_i <= 3'b010;    //+
			7'd10: rom_i <= 3'b110;   //[
			7'd11: rom_i <= 3'b001;   //>
			7'd12: rom_i <= 3'b010;   //+
			7'd13: rom_i <= 3'b010;   //+
			7'd14: rom_i <= 3'b010;   //+
			7'd15: rom_i <= 3'b010;   //+
			7'd16: rom_i <= 3'b010;   //+
			7'd17: rom_i <= 3'b010;   //+
			7'd18: rom_i <= 3'b010;   //+
			7'd19: rom_i <= 3'b001;   //>
			7'd20: rom_i <= 3'b010;   //+
			7'd21: rom_i <= 3'b010;   //+
			7'd22: rom_i <= 3'b010;   //+
			7'd23: rom_i <= 3'b010;   //+
			7'd24: rom_i <= 3'b010;   //+
			7'd25: rom_i <= 3'b010;   //+
			7'd26: rom_i <= 3'b010;   //+
			7'd27: rom_i <= 3'b010;   //+
			7'd28: rom_i <= 3'b010;   //+
			7'd29: rom_i <= 3'b010;   //+
			7'd30: rom_i <= 3'b001;   //>
			7'd31: rom_i <= 3'b010;   //+
			7'd32: rom_i <= 3'b010;   //+
			7'd33: rom_i <= 3'b010;   //+
			7'd34: rom_i <= 3'b001;   //>
			7'd35: rom_i <= 3'b010;   //+
			7'd36: rom_i <= 3'b000;   //<
			7'd37: rom_i <= 3'b000;   //<
			7'd38: rom_i <= 3'b000;   //<
			7'd39: rom_i <= 3'b000;   //<
			7'd40: rom_i <= 3'b011;   //-
			7'd41: rom_i <= 3'b111;   //]
			7'd42: rom_i <= 3'b001;   //>
			7'd43: rom_i <= 3'b010;   //+
			7'd44: rom_i <= 3'b010;   //+
			7'd45: rom_i <= 3'b101;   //.
			7'd46: rom_i <= 3'b001;   //>
			7'd47: rom_i <= 3'b010;   //+
			7'd48: rom_i <= 3'b101;   //.
			7'd49: rom_i <= 3'b010;   //+
			7'd50: rom_i <= 3'b010;   //+
			7'd51: rom_i <= 3'b010;   //+
			7'd52: rom_i <= 3'b010;   //+
			7'd53: rom_i <= 3'b010;   //+
			7'd54: rom_i <= 3'b010;   //+
			7'd55: rom_i <= 3'b010;   //+
			7'd56: rom_i <= 3'b101;   //.
			7'd57: rom_i <= 3'b101;   //.
			7'd58: rom_i <= 3'b010;   //+
			7'd59: rom_i <= 3'b010;   //+
			7'd60: rom_i <= 3'b010;   //+
			7'd61: rom_i <= 3'b101;   //.
			7'd62: rom_i <= 3'b001;   //>
			7'd63: rom_i <= 3'b010;   //+
			7'd64: rom_i <= 3'b010;   //+
			7'd65: rom_i <= 3'b101;   //.
			7'd66: rom_i <= 3'b000;   //<
			7'd67: rom_i <= 3'b000;   //<
			7'd68: rom_i <= 3'b010;   //+
			7'd69: rom_i <= 3'b010;   //+
			7'd70: rom_i <= 3'b010;   //+
			7'd71: rom_i <= 3'b010;   //+
			7'd72: rom_i <= 3'b010;   //+
			7'd73: rom_i <= 3'b010;   //+
			7'd74: rom_i <= 3'b010;   //+
			7'd75: rom_i <= 3'b010;   //+
			7'd76: rom_i <= 3'b010;   //+
			7'd77: rom_i <= 3'b010;   //+
			7'd78: rom_i <= 3'b010;   //+
			7'd79: rom_i <= 3'b010;   //+
			7'd80: rom_i <= 3'b010;   //+
			7'd81: rom_i <= 3'b010;   //+
			7'd82: rom_i <= 3'b010;   //+
			7'd83: rom_i <= 3'b101;   //.
			7'd84: rom_i <= 3'b001;   //>
			7'd85: rom_i <= 3'b101;   //.
			7'd86: rom_i <= 3'b010;   //+
			7'd87: rom_i <= 3'b010;   //+
			7'd88: rom_i <= 3'b010;   //+
			7'd89: rom_i <= 3'b101;   //.
			7'd90: rom_i <= 3'b011;   //-
			7'd91: rom_i <= 3'b011;   //-
			7'd92: rom_i <= 3'b011;   //-
			7'd93: rom_i <= 3'b011;   //-
			7'd94: rom_i <= 3'b011;   //-
			7'd95: rom_i <= 3'b011;   //-
			7'd96: rom_i <= 3'b101;   //.
			7'd97: rom_i <= 3'b011;   //-
			7'd98: rom_i <= 3'b011;   //-
			7'd99: rom_i <= 3'b011;   //-
			7'd100: rom_i <= 3'b011;  //-
			7'd101: rom_i <= 3'b011;  //-
			7'd102: rom_i <= 3'b011;  //-
			7'd103: rom_i <= 3'b011;  //-
			7'd104: rom_i <= 3'b011;  //-
			7'd105: rom_i <= 3'b101;  //.
			7'd106: rom_i <= 3'b001;  //>
			7'd107: rom_i <= 3'b010;  //+
			7'd108: rom_i <= 3'b101;  //.
			7'd109: rom_i <= 3'b001;  //>
			7'd110: rom_i <= 3'b101;  //.
			7'd111: rom_i <= 3'b110;  //[
			7'd112: rom_i <= 3'b010;  //+
			7'd113: rom_i <= 3'b011;  //-
			7'd114: rom_i <= 3'b111;  //]
			7'd115: rom_i <= 3'b000;
			7'd116: rom_i <= 3'b000;
			7'd117: rom_i <= 3'b000;
			7'd118: rom_i <= 3'b000;
			7'd119: rom_i <= 3'b000;
			7'd120: rom_i <= 3'b000;
			7'd121: rom_i <= 3'b000;
			7'd122: rom_i <= 3'b000;
			7'd123: rom_i <= 3'b000;
			7'd124: rom_i <= 3'b000;
			7'd125: rom_i <= 3'b000;
			7'd126: rom_i <= 3'b000;
			7'd127: rom_i <= 3'b000;

		endcase
	end

endmodule
